`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: Ashot Hambardzumyan
// 
// Create Date: 10/27/2016 05:57:13 PM
// Design Name: 
// Module Name: road
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module road(
input wire clk, reset,refresh_tick, pause,enter_key,
input wire [9:0] pixel_x, pixel_y,
output wire road_on, output reg finish_line, //i can add output obstacle_x as a line or two pixels on the road, they will be red
output reg [11:0] road_rgb,
output reg [11:0] obstacle_rgb
);

//variables 
//square canvas for the road 




localparam MAX_X = 512;
localparam MAX_Y = 480;
localparam road_x_l = 64;
localparam road_x_r = road_x_l + MAX_X-1;
localparam road_y_t = 0;
localparam road_y_b = MAX_Y-1;
localparam road_x_delta = 120; //thickness of the road
 
reg [9:0] road_rom_addr; //960 lines
reg [8:0] road_rom_col; //512 lines
reg [0:511] road_rom_data; //x data length
wire road_rom_bit, canvas_on;
reg [11:0] counter, tempC;
reg [1:0] finish;
reg slow_count; //[1:0]

//adding obstacle

//reg[9:0] obstacle_x;


assign canvas_on =  (road_x_l<=pixel_x) && (pixel_x<=road_x_r);
assign road_rom_bit = road_rom_data[road_rom_col];
assign road_on = canvas_on & road_rom_bit;

//rolling road
always@(posedge clk)
begin
if(reset)
    begin
    // reset the road position,
    // sets the road such that car is at a flat part of the road
    counter <=4*MAX_Y -440; 
    finish <= 0;
    end
//if paused, don't increament the counter, pause the movement
else if(refresh_tick && !pause) 
    begin
     counter <= tempC%(4*MAX_Y);
     if((counter !=44)&& 
     (tempC%(4*MAX_Y) == 42 || tempC%(4*MAX_Y) == 44)) 
           finish <= finish + 1;
    end
else
    begin // this part could have been in else if.
    //it is here because gate level path was too long 
    if(enter_key) //turbo, road moves 2X the speed
     tempC <= (counter + 4*MAX_Y - 4);
    else
     tempC <= (counter + 4*MAX_Y - 2);
    end

    
//making this a reg so that synthesiser inferes ram
road_rom_addr <= (pixel_y + counter)%(2*MAX_Y);


//indexing scheme: I use the original 2 frames 
//for frame 3 and 4, by fliping 1, 2 from left to right
//for a data that is power of 2, fliping LR is simple
//just invert the bit index
if(((pixel_y + counter)%(4*MAX_Y))>(2*MAX_Y))
   begin
   road_rom_col <= ~(pixel_x[8:0]-road_x_l);
   end
else
   begin
   road_rom_col <= (pixel_x[8:0]-road_x_l);
   end
  
end


always@*
begin
//wait for 8 frames, before enabling finish line, 
  //show the finish line
  if(road_rom_addr == 0 && (finish==2))
      begin;
        finish_line =1'b1;
        road_rgb = 12'hf00;
      end
// wait for 4 frames i guess before having an obstacle or just add it in initial frames
// else if(road_rom_addr==0 && (finish==0))
//        begin
//          road_rgb=12'hff0; // this adds a yellow line which can act as point
          
//      end
      else
          begin
           obstacle_rgb=12'hff0;
           road_rgb = 12'h555; //changes
           finish_line = 1'b0;
          end
  

end

//960 lines of bitmap for the road. 2 full frames at 480 lines per frame.
// using indexing scheme above the 2 frames become 4 frames, that roll continuesly
//looping back to itself.
//Below is the C# code for generating this road. I used 2 sine waves, 
// to genearte this road.
/*
static void Main(string[] args)
        {
        int[] ver = new int[960];
        for (int i = 0; i < 960; i++)
        {
                if (i < 50)
                    ver[i] = 256;
                else if (i < 910)
                    ver[i] = (int)Math.Floor(-256 * 0.5 * (Math.Sin((i - 50) * Math.PI / 430)
                        + 0.75 * Math.Sin((i - 50) * 0.5 * Math.PI / 430))) + 256;
                else
                    ver[i] = 256;
                if (ver[i] <100)
                {
                ver[i] = 100;
                }
                else if (ver[i] > 412)
                {
                    ver[i] = 412;
                }
        }
        String temp = null;
        for (int i = 0; i < 960; i++)
        {
            //9'd000: road_rom_data = {220'b0,{72{1'b1}},220'b0}; 
            temp = "10'd" + i + ": road_rom_data = {" + (ver[i]-60)+ "'b0,{"
                    + 120 + "{1'b1}}," + (512 - 60 - ver[i]) + "'b0};";
                Console.WriteLine(temp);
        }
    }

*/


always @*
  case(road_rom_addr)
  10'd0: road_rom_data = {220'b0,{72{1'b1}},220'b0};
  10'd1: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd2: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd3: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd4: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd5: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd6: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd7: road_rom_data = {220'b0,{96{1'b1}},196'b0};
  10'd8: road_rom_data = {220'b0,{96{1'b1}},196'b0};
  10'd9: road_rom_data = {220'b0,{96{1'b1}},196'b0};
  10'd10: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd11: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd12: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd13: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd14: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd15: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd16: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd17: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd18: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd19: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd20: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd21: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd22: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd23: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd24: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd25: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd26: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd27: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd28: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd29: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd30: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd31: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd32: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd33: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd34: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd35: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd36: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd37: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd38: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd39: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd40: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd41: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd42: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd43: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd44: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd45: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd46: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd47: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd48: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd49: road_rom_data = {200'b0,{114{1'b1}},198'b0};//bringing in obstacle green
  10'd50: road_rom_data = {200'b0,{114{1'b1}},198'b0};//bringing in obstacle green
  10'd51: road_rom_data = {200'b0,{114{1'b1}},198'b0};//bringing in obstacle green
  10'd52: road_rom_data = {193'b0,{120{1'b1}},199'b0};
  10'd53: road_rom_data = {192'b0,{120{1'b1}},200'b0};
  10'd54: road_rom_data = {190'b0,{120{1'b1}},202'b0};
  10'd55: road_rom_data = {189'b0,{120{1'b1}},203'b0};
  10'd56: road_rom_data = {188'b0,{120{1'b1}},204'b0};
  10'd57: road_rom_data = {187'b0,{120{1'b1}},205'b0};
  10'd58: road_rom_data = {185'b0,{120{1'b1}},207'b0};
  10'd59: road_rom_data = {184'b0,{120{1'b1}},208'b0};
  10'd60: road_rom_data = {183'b0,{120{1'b1}},209'b0};
  10'd61: road_rom_data = {181'b0,{120{1'b1}},211'b0};
  10'd62: road_rom_data = {180'b0,{120{1'b1}},212'b0};
  10'd63: road_rom_data = {179'b0,{120{1'b1}},213'b0};
  10'd64: road_rom_data = {178'b0,{120{1'b1}},214'b0};
  10'd65: road_rom_data = {176'b0,{120{1'b1}},216'b0};
  10'd66: road_rom_data = {175'b0,{120{1'b1}},217'b0};
  10'd67: road_rom_data = {174'b0,{120{1'b1}},218'b0};
  10'd68: road_rom_data = {172'b0,{120{1'b1}},220'b0};
  10'd69: road_rom_data = {171'b0,{120{1'b1}},221'b0};
  10'd70: road_rom_data = {170'b0,{120{1'b1}},222'b0};
  10'd71: road_rom_data = {169'b0,{120{1'b1}},223'b0};
  10'd72: road_rom_data = {167'b0,{120{1'b1}},225'b0};
  10'd73: road_rom_data = {166'b0,{120{1'b1}},226'b0};
  10'd74: road_rom_data = {165'b0,{120{1'b1}},227'b0};
  10'd75: road_rom_data = {163'b0,{120{1'b1}},229'b0};
  10'd76: road_rom_data = {162'b0,{120{1'b1}},230'b0};
  10'd77: road_rom_data = {161'b0,{120{1'b1}},231'b0};
  10'd78: road_rom_data = {160'b0,{120{1'b1}},232'b0};
  10'd79: road_rom_data = {158'b0,{120{1'b1}},234'b0};
  10'd80: road_rom_data = {157'b0,{120{1'b1}},235'b0};
  10'd81: road_rom_data = {156'b0,{120{1'b1}},236'b0};
  10'd82: road_rom_data = {155'b0,{120{1'b1}},237'b0};
  10'd83: road_rom_data = {153'b0,{120{1'b1}},239'b0};
  10'd84: road_rom_data = {152'b0,{120{1'b1}},240'b0};
  10'd85: road_rom_data = {151'b0,{120{1'b1}},241'b0};
  10'd86: road_rom_data = {150'b0,{120{1'b1}},242'b0};
  10'd87: road_rom_data = {148'b0,{120{1'b1}},244'b0};
  10'd88: road_rom_data = {147'b0,{120{1'b1}},245'b0};
  10'd89: road_rom_data = {146'b0,{120{1'b1}},246'b0};
  10'd90: road_rom_data = {145'b0,{120{1'b1}},247'b0};
  10'd91: road_rom_data = {143'b0,{120{1'b1}},249'b0};
  10'd92: road_rom_data = {142'b0,{120{1'b1}},250'b0};
  10'd93: road_rom_data = {141'b0,{120{1'b1}},251'b0};
  10'd94: road_rom_data = {140'b0,{120{1'b1}},252'b0};
  10'd95: road_rom_data = {138'b0,{120{1'b1}},254'b0};
  10'd96: road_rom_data = {137'b0,{120{1'b1}},255'b0};
  10'd97: road_rom_data = {136'b0,{120{1'b1}},256'b0};
  10'd98: road_rom_data = {135'b0,{120{1'b1}},257'b0};
  10'd99: road_rom_data = {134'b0,{120{1'b1}},258'b0};
  10'd100: road_rom_data = {132'b0,{120{1'b1}},260'b0};
  10'd101: road_rom_data = {131'b0,{120{1'b1}},261'b0};
  10'd102: road_rom_data = {130'b0,{120{1'b1}},262'b0};
  10'd103: road_rom_data = {129'b0,{120{1'b1}},263'b0};
  10'd104: road_rom_data = {127'b0,{120{1'b1}},265'b0};
  10'd105: road_rom_data = {126'b0,{120{1'b1}},266'b0};
  10'd106: road_rom_data = {125'b0,{120{1'b1}},267'b0};
  10'd107: road_rom_data = {124'b0,{120{1'b1}},268'b0};
  10'd108: road_rom_data = {123'b0,{120{1'b1}},269'b0};
  10'd109: road_rom_data = {121'b0,{120{1'b1}},271'b0};
  10'd110: road_rom_data = {120'b0,{120{1'b1}},272'b0};
  10'd111: road_rom_data = {119'b0,{120{1'b1}},273'b0};
  10'd112: road_rom_data = {118'b0,{120{1'b1}},274'b0};
  10'd113: road_rom_data = {117'b0,{120{1'b1}},275'b0};
  10'd114: road_rom_data = {116'b0,{120{1'b1}},276'b0};
  10'd115: road_rom_data = {114'b0,{120{1'b1}},278'b0};
  10'd116: road_rom_data = {113'b0,{120{1'b1}},279'b0};
  10'd117: road_rom_data = {112'b0,{120{1'b1}},280'b0};
  10'd118: road_rom_data = {111'b0,{120{1'b1}},281'b0};
  10'd119: road_rom_data = {110'b0,{120{1'b1}},282'b0};
  10'd120: road_rom_data = {109'b0,{120{1'b1}},283'b0};
  10'd121: road_rom_data = {107'b0,{120{1'b1}},285'b0};
  10'd122: road_rom_data = {106'b0,{120{1'b1}},286'b0};
  10'd123: road_rom_data = {105'b0,{120{1'b1}},287'b0};
  10'd124: road_rom_data = {104'b0,{120{1'b1}},288'b0};
  10'd125: road_rom_data = {103'b0,{120{1'b1}},289'b0};
  10'd126: road_rom_data = {102'b0,{120{1'b1}},290'b0};
  10'd127: road_rom_data = {101'b0,{120{1'b1}},291'b0};
  10'd128: road_rom_data = {99'b0,{120{1'b1}},293'b0};
  10'd129: road_rom_data = {98'b0,{120{1'b1}},294'b0};
  10'd130: road_rom_data = {97'b0,{120{1'b1}},295'b0};
  10'd131: road_rom_data = {96'b0,{120{1'b1}},296'b0};
  10'd132: road_rom_data = {95'b0,{120{1'b1}},297'b0};
  10'd133: road_rom_data = {94'b0,{120{1'b1}},298'b0};
  10'd134: road_rom_data = {93'b0,{120{1'b1}},299'b0};
  10'd135: road_rom_data = {92'b0,{120{1'b1}},300'b0};
  10'd136: road_rom_data = {91'b0,{120{1'b1}},301'b0};
  10'd137: road_rom_data = {90'b0,{120{1'b1}},302'b0};
  10'd138: road_rom_data = {88'b0,{120{1'b1}},304'b0};
  10'd139: road_rom_data = {87'b0,{120{1'b1}},305'b0};
  10'd140: road_rom_data = {86'b0,{120{1'b1}},306'b0};
  10'd141: road_rom_data = {85'b0,{120{1'b1}},307'b0};
  10'd142: road_rom_data = {84'b0,{120{1'b1}},308'b0};
  10'd143: road_rom_data = {83'b0,{120{1'b1}},309'b0};
  10'd144: road_rom_data = {82'b0,{120{1'b1}},310'b0};
  10'd145: road_rom_data = {81'b0,{120{1'b1}},311'b0};
  10'd146: road_rom_data = {80'b0,{120{1'b1}},312'b0};
  10'd147: road_rom_data = {79'b0,{120{1'b1}},313'b0};
  10'd148: road_rom_data = {78'b0,{120{1'b1}},314'b0};
  10'd149: road_rom_data = {77'b0,{120{1'b1}},315'b0};
  10'd150: road_rom_data = {76'b0,{120{1'b1}},316'b0};
  10'd151: road_rom_data = {75'b0,{120{1'b1}},317'b0};
  10'd152: road_rom_data = {74'b0,{120{1'b1}},318'b0};
  10'd153: road_rom_data = {73'b0,{120{1'b1}},319'b0};
  10'd154: road_rom_data = {72'b0,{120{1'b1}},320'b0};
  10'd155: road_rom_data = {71'b0,{120{1'b1}},321'b0};
  10'd156: road_rom_data = {70'b0,{120{1'b1}},322'b0};
  10'd157: road_rom_data = {69'b0,{120{1'b1}},323'b0};
  10'd158: road_rom_data = {68'b0,{120{1'b1}},324'b0};
  10'd159: road_rom_data = {67'b0,{120{1'b1}},325'b0};
  10'd160: road_rom_data = {66'b0,{120{1'b1}},326'b0};
  10'd161: road_rom_data = {65'b0,{120{1'b1}},327'b0};
  10'd162: road_rom_data = {64'b0,{120{1'b1}},328'b0};
  10'd163: road_rom_data = {63'b0,{120{1'b1}},329'b0};
  10'd164: road_rom_data = {62'b0,{120{1'b1}},330'b0};
  10'd165: road_rom_data = {61'b0,{120{1'b1}},331'b0};
  10'd166: road_rom_data = {60'b0,{120{1'b1}},332'b0};
  10'd167: road_rom_data = {59'b0,{120{1'b1}},333'b0};
  10'd168: road_rom_data = {58'b0,{120{1'b1}},334'b0};
  10'd169: road_rom_data = {57'b0,{120{1'b1}},335'b0};
  10'd170: road_rom_data = {56'b0,{120{1'b1}},336'b0};
  10'd171: road_rom_data = {55'b0,{120{1'b1}},337'b0};
  10'd172: road_rom_data = {55'b0,{120{1'b1}},337'b0};
  10'd173: road_rom_data = {54'b0,{120{1'b1}},338'b0};
  10'd174: road_rom_data = {53'b0,{120{1'b1}},339'b0};
  10'd175: road_rom_data = {52'b0,{120{1'b1}},340'b0};
  10'd176: road_rom_data = {51'b0,{120{1'b1}},341'b0};
  10'd177: road_rom_data = {50'b0,{120{1'b1}},342'b0};
  10'd178: road_rom_data = {49'b0,{120{1'b1}},343'b0};
  10'd179: road_rom_data = {48'b0,{120{1'b1}},344'b0};
  10'd180: road_rom_data = {48'b0,{120{1'b1}},344'b0};
  10'd181: road_rom_data = {47'b0,{120{1'b1}},345'b0};
  10'd182: road_rom_data = {46'b0,{120{1'b1}},346'b0};
  10'd183: road_rom_data = {45'b0,{120{1'b1}},347'b0};
  10'd184: road_rom_data = {44'b0,{120{1'b1}},348'b0};
  10'd185: road_rom_data = {43'b0,{120{1'b1}},349'b0};
  10'd186: road_rom_data = {42'b0,{120{1'b1}},350'b0};
  10'd187: road_rom_data = {42'b0,{120{1'b1}},350'b0};
  10'd188: road_rom_data = {41'b0,{120{1'b1}},351'b0};
  10'd189: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd190: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd191: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd192: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd193: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd194: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd195: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd196: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd197: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd198: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd199: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd200: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd201: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd202: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd203: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd204: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd205: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd206: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd207: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd208: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd209: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd210: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd211: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd212: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd213: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd214: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd215: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd216: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd217: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd218: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd219: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd220: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd221: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd222: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd223: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd224: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd225: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd226: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd227: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd228: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd229: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd230: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd231: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd232: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd233: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd234: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd235: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd236: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd237: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd238: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd239: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd240: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd241: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd242: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd243: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd244: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd245: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd246: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd247: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd248: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd249: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd250: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd251: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd252: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd253: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd254: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd255: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd256: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd257: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd258: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd259: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd260: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd261: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd262: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd263: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd264: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd265: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd266: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd267: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd268: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd269: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd270: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd271: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd272: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd273: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd274: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd275: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd276: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd277: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd278: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd279: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd280: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd281: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd282: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd283: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd284: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd285: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd286: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd287: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd288: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd289: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd290: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd291: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd292: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd293: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd294: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd295: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd296: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd297: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd298: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd299: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd300: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd301: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd302: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd303: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd304: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd305: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd306: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd307: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd308: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd309: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd310: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd311: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd312: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd313: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd314: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd315: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd316: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd317: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd318: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd319: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd320: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd321: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd322: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd323: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd324: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd325: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd326: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd327: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd328: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd329: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd330: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd331: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd332: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd333: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd334: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd335: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd336: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd337: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd338: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd339: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd340: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd341: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd342: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd343: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd344: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd345: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd346: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd347: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd348: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd349: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd350: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd351: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd352: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd353: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd354: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd355: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd356: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd357: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd358: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd359: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd360: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd361: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd362: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd363: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd364: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd365: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd366: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd367: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd368: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd369: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd370: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd371: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd372: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd373: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd374: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd375: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd376: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd377: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd378: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd379: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd380: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd381: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd382: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd383: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd384: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd385: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd386: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd387: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd388: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd389: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd390: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd391: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd392: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd393: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd394: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd395: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd396: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd397: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd398: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd399: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd400: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd401: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd402: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd403: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd404: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd405: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd406: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd407: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd408: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd409: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd410: road_rom_data = {40'b0,{120{1'b1}},352'b0};
  10'd411: road_rom_data = {41'b0,{120{1'b1}},351'b0};
  10'd412: road_rom_data = {41'b0,{120{1'b1}},351'b0};
  10'd413: road_rom_data = {42'b0,{120{1'b1}},350'b0};
  10'd414: road_rom_data = {43'b0,{120{1'b1}},349'b0};
  10'd415: road_rom_data = {44'b0,{120{1'b1}},348'b0};
  10'd416: road_rom_data = {44'b0,{120{1'b1}},348'b0};
  10'd417: road_rom_data = {45'b0,{120{1'b1}},347'b0};
  10'd418: road_rom_data = {46'b0,{120{1'b1}},346'b0};
  10'd419: road_rom_data = {47'b0,{120{1'b1}},345'b0};
  10'd420: road_rom_data = {47'b0,{120{1'b1}},345'b0};
  10'd421: road_rom_data = {48'b0,{120{1'b1}},344'b0};
  10'd422: road_rom_data = {49'b0,{120{1'b1}},343'b0};
  10'd423: road_rom_data = {50'b0,{120{1'b1}},342'b0};
  10'd424: road_rom_data = {51'b0,{120{1'b1}},341'b0};
  10'd425: road_rom_data = {51'b0,{120{1'b1}},341'b0};
  10'd426: road_rom_data = {52'b0,{120{1'b1}},340'b0};
  10'd427: road_rom_data = {53'b0,{120{1'b1}},339'b0};
  10'd428: road_rom_data = {54'b0,{120{1'b1}},338'b0};
  10'd429: road_rom_data = {55'b0,{120{1'b1}},337'b0};
  10'd430: road_rom_data = {55'b0,{120{1'b1}},337'b0};
  10'd431: road_rom_data = {56'b0,{120{1'b1}},336'b0};
  10'd432: road_rom_data = {57'b0,{120{1'b1}},335'b0};
  10'd433: road_rom_data = {58'b0,{120{1'b1}},334'b0};
  10'd434: road_rom_data = {59'b0,{120{1'b1}},333'b0};
  10'd435: road_rom_data = {59'b0,{120{1'b1}},333'b0};
  10'd436: road_rom_data = {60'b0,{120{1'b1}},332'b0};
  10'd437: road_rom_data = {61'b0,{120{1'b1}},331'b0};
  10'd438: road_rom_data = {62'b0,{120{1'b1}},330'b0};
  10'd439: road_rom_data = {63'b0,{120{1'b1}},329'b0};
  10'd440: road_rom_data = {64'b0,{120{1'b1}},328'b0};
  10'd441: road_rom_data = {64'b0,{120{1'b1}},328'b0};
  10'd442: road_rom_data = {65'b0,{120{1'b1}},327'b0};
  10'd443: road_rom_data = {66'b0,{120{1'b1}},326'b0};
  10'd444: road_rom_data = {67'b0,{120{1'b1}},325'b0};
  10'd445: road_rom_data = {68'b0,{120{1'b1}},324'b0};
  10'd446: road_rom_data = {69'b0,{120{1'b1}},323'b0};
  10'd447: road_rom_data = {70'b0,{120{1'b1}},322'b0};
  10'd448: road_rom_data = {71'b0,{120{1'b1}},321'b0};
  10'd449: road_rom_data = {71'b0,{120{1'b1}},321'b0};
  10'd450: road_rom_data = {72'b0,{120{1'b1}},320'b0};
  10'd451: road_rom_data = {73'b0,{120{1'b1}},319'b0};
  10'd452: road_rom_data = {74'b0,{120{1'b1}},318'b0};
  10'd453: road_rom_data = {75'b0,{120{1'b1}},317'b0};
  10'd454: road_rom_data = {76'b0,{120{1'b1}},316'b0};
  10'd455: road_rom_data = {77'b0,{120{1'b1}},315'b0};
  10'd456: road_rom_data = {78'b0,{120{1'b1}},314'b0};
  10'd457: road_rom_data = {78'b0,{120{1'b1}},314'b0};
  10'd458: road_rom_data = {79'b0,{120{1'b1}},313'b0};
  10'd459: road_rom_data = {80'b0,{120{1'b1}},312'b0};
  10'd460: road_rom_data = {81'b0,{120{1'b1}},311'b0};
  10'd461: road_rom_data = {82'b0,{120{1'b1}},310'b0};
  10'd462: road_rom_data = {83'b0,{120{1'b1}},309'b0};
  10'd463: road_rom_data = {84'b0,{120{1'b1}},308'b0};
  10'd464: road_rom_data = {85'b0,{120{1'b1}},307'b0};
  10'd465: road_rom_data = {86'b0,{120{1'b1}},306'b0};
  10'd466: road_rom_data = {87'b0,{120{1'b1}},305'b0};
  10'd467: road_rom_data = {87'b0,{120{1'b1}},305'b0};
  10'd468: road_rom_data = {88'b0,{120{1'b1}},304'b0};
  10'd469: road_rom_data = {89'b0,{120{1'b1}},303'b0};
  10'd470: road_rom_data = {90'b0,{120{1'b1}},302'b0};
  10'd471: road_rom_data = {91'b0,{120{1'b1}},301'b0};
  10'd472: road_rom_data = {92'b0,{120{1'b1}},300'b0};
  10'd473: road_rom_data = {93'b0,{120{1'b1}},299'b0};
  10'd474: road_rom_data = {94'b0,{120{1'b1}},298'b0};
  10'd475: road_rom_data = {95'b0,{120{1'b1}},297'b0};
  10'd476: road_rom_data = {96'b0,{120{1'b1}},296'b0};
  10'd477: road_rom_data = {97'b0,{120{1'b1}},295'b0};
  10'd478: road_rom_data = {98'b0,{120{1'b1}},294'b0};
  10'd479: road_rom_data = {99'b0,{120{1'b1}},293'b0};
  10'd480: road_rom_data = {99'b0,{120{1'b1}},293'b0};
  10'd481: road_rom_data = {100'b0,{120{1'b1}},292'b0};
  10'd482: road_rom_data = {101'b0,{120{1'b1}},291'b0};
  10'd483: road_rom_data = {102'b0,{120{1'b1}},290'b0};
  10'd484: road_rom_data = {103'b0,{120{1'b1}},289'b0};
  10'd485: road_rom_data = {104'b0,{120{1'b1}},288'b0};
  10'd486: road_rom_data = {105'b0,{120{1'b1}},287'b0};
  10'd487: road_rom_data = {106'b0,{120{1'b1}},286'b0};
  10'd488: road_rom_data = {107'b0,{120{1'b1}},285'b0};
  10'd489: road_rom_data = {108'b0,{120{1'b1}},284'b0};
  10'd490: road_rom_data = {109'b0,{120{1'b1}},283'b0};
  10'd491: road_rom_data = {110'b0,{120{1'b1}},282'b0};
  10'd492: road_rom_data = {111'b0,{120{1'b1}},281'b0};
  10'd493: road_rom_data = {112'b0,{120{1'b1}},280'b0};
  10'd494: road_rom_data = {113'b0,{120{1'b1}},279'b0};
  10'd495: road_rom_data = {114'b0,{120{1'b1}},278'b0};
  10'd496: road_rom_data = {115'b0,{120{1'b1}},277'b0};
  10'd497: road_rom_data = {116'b0,{120{1'b1}},276'b0};
  10'd498: road_rom_data = {116'b0,{120{1'b1}},276'b0};
  10'd499: road_rom_data = {117'b0,{120{1'b1}},275'b0};
  10'd500: road_rom_data = {118'b0,{120{1'b1}},274'b0};
  10'd501: road_rom_data = {119'b0,{120{1'b1}},273'b0};
  10'd502: road_rom_data = {120'b0,{120{1'b1}},272'b0};
  10'd503: road_rom_data = {121'b0,{120{1'b1}},271'b0};
  10'd504: road_rom_data = {122'b0,{120{1'b1}},270'b0};
  10'd505: road_rom_data = {123'b0,{120{1'b1}},269'b0};
  10'd506: road_rom_data = {124'b0,{120{1'b1}},268'b0};
  10'd507: road_rom_data = {125'b0,{120{1'b1}},267'b0};
  10'd508: road_rom_data = {126'b0,{120{1'b1}},266'b0};
  10'd509: road_rom_data = {127'b0,{120{1'b1}},265'b0};
  10'd510: road_rom_data = {128'b0,{120{1'b1}},264'b0};
  10'd511: road_rom_data = {129'b0,{120{1'b1}},263'b0};
  10'd512: road_rom_data = {130'b0,{120{1'b1}},262'b0};
  10'd513: road_rom_data = {131'b0,{120{1'b1}},261'b0};
  10'd514: road_rom_data = {132'b0,{120{1'b1}},260'b0};
  10'd515: road_rom_data = {133'b0,{120{1'b1}},259'b0};
  10'd516: road_rom_data = {134'b0,{120{1'b1}},258'b0};
  10'd517: road_rom_data = {135'b0,{120{1'b1}},257'b0};
  10'd518: road_rom_data = {136'b0,{120{1'b1}},256'b0};
  10'd519: road_rom_data = {136'b0,{120{1'b1}},256'b0};
  10'd520: road_rom_data = {137'b0,{120{1'b1}},255'b0};
  10'd521: road_rom_data = {138'b0,{120{1'b1}},254'b0};
  10'd522: road_rom_data = {139'b0,{120{1'b1}},253'b0};
  10'd523: road_rom_data = {140'b0,{120{1'b1}},252'b0};
  10'd524: road_rom_data = {141'b0,{120{1'b1}},251'b0};
  10'd525: road_rom_data = {142'b0,{120{1'b1}},250'b0};
  10'd526: road_rom_data = {143'b0,{120{1'b1}},249'b0};
  10'd527: road_rom_data = {144'b0,{120{1'b1}},248'b0};
  10'd528: road_rom_data = {145'b0,{120{1'b1}},247'b0};
  10'd529: road_rom_data = {146'b0,{120{1'b1}},246'b0};
  10'd530: road_rom_data = {147'b0,{120{1'b1}},245'b0};
  10'd531: road_rom_data = {148'b0,{120{1'b1}},244'b0};
  10'd532: road_rom_data = {149'b0,{120{1'b1}},243'b0};
  10'd533: road_rom_data = {150'b0,{120{1'b1}},242'b0};
  10'd534: road_rom_data = {151'b0,{120{1'b1}},241'b0};
  10'd535: road_rom_data = {151'b0,{120{1'b1}},241'b0};
  10'd536: road_rom_data = {152'b0,{120{1'b1}},240'b0};
  10'd537: road_rom_data = {153'b0,{120{1'b1}},239'b0};
  10'd538: road_rom_data = {154'b0,{120{1'b1}},238'b0};
  10'd539: road_rom_data = {155'b0,{120{1'b1}},237'b0};
  10'd540: road_rom_data = {156'b0,{120{1'b1}},236'b0};
  10'd541: road_rom_data = {157'b0,{120{1'b1}},235'b0};
  10'd542: road_rom_data = {158'b0,{120{1'b1}},234'b0};
  10'd543: road_rom_data = {159'b0,{120{1'b1}},233'b0};
  10'd544: road_rom_data = {160'b0,{120{1'b1}},232'b0};
  10'd545: road_rom_data = {161'b0,{120{1'b1}},231'b0};
  10'd546: road_rom_data = {162'b0,{120{1'b1}},230'b0};
  10'd547: road_rom_data = {163'b0,{120{1'b1}},229'b0};
  10'd548: road_rom_data = {163'b0,{120{1'b1}},229'b0};
  10'd549: road_rom_data = {164'b0,{120{1'b1}},228'b0};
  10'd550: road_rom_data = {165'b0,{120{1'b1}},227'b0};
  10'd551: road_rom_data = {166'b0,{120{1'b1}},226'b0};
  10'd552: road_rom_data = {167'b0,{120{1'b1}},225'b0};
  10'd553: road_rom_data = {168'b0,{120{1'b1}},224'b0};
  10'd554: road_rom_data = {169'b0,{120{1'b1}},223'b0};
  10'd555: road_rom_data = {170'b0,{120{1'b1}},222'b0};
  10'd556: road_rom_data = {171'b0,{120{1'b1}},221'b0};
  10'd557: road_rom_data = {172'b0,{120{1'b1}},220'b0};
  10'd558: road_rom_data = {172'b0,{120{1'b1}},220'b0};
  10'd559: road_rom_data = {173'b0,{120{1'b1}},219'b0};
  10'd560: road_rom_data = {174'b0,{120{1'b1}},218'b0};
  10'd561: road_rom_data = {175'b0,{120{1'b1}},217'b0};
  10'd562: road_rom_data = {176'b0,{120{1'b1}},216'b0};
  10'd563: road_rom_data = {177'b0,{120{1'b1}},215'b0};
  10'd564: road_rom_data = {178'b0,{120{1'b1}},214'b0};
  10'd565: road_rom_data = {179'b0,{120{1'b1}},213'b0};
  10'd566: road_rom_data = {179'b0,{120{1'b1}},213'b0};
  10'd567: road_rom_data = {180'b0,{120{1'b1}},212'b0};
  10'd568: road_rom_data = {181'b0,{120{1'b1}},211'b0};
  10'd569: road_rom_data = {182'b0,{120{1'b1}},210'b0};
  10'd570: road_rom_data = {183'b0,{120{1'b1}},209'b0};
  10'd571: road_rom_data = {184'b0,{120{1'b1}},208'b0};
  10'd572: road_rom_data = {185'b0,{120{1'b1}},207'b0};
  10'd573: road_rom_data = {185'b0,{120{1'b1}},207'b0};
  10'd574: road_rom_data = {186'b0,{120{1'b1}},206'b0};
  10'd575: road_rom_data = {187'b0,{120{1'b1}},205'b0};
  10'd576: road_rom_data = {188'b0,{120{1'b1}},204'b0};
  10'd577: road_rom_data = {189'b0,{120{1'b1}},203'b0};
  10'd578: road_rom_data = {190'b0,{120{1'b1}},202'b0};
  10'd579: road_rom_data = {190'b0,{120{1'b1}},202'b0};
  10'd580: road_rom_data = {191'b0,{120{1'b1}},201'b0};
  10'd581: road_rom_data = {192'b0,{120{1'b1}},200'b0};
  10'd582: road_rom_data = {193'b0,{120{1'b1}},199'b0};
  10'd583: road_rom_data = {194'b0,{120{1'b1}},198'b0};
  10'd584: road_rom_data = {195'b0,{120{1'b1}},197'b0};
  10'd585: road_rom_data = {195'b0,{120{1'b1}},197'b0};
  10'd586: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd587: road_rom_data = {197'b0,{120{1'b1}},195'b0};
  10'd588: road_rom_data = {198'b0,{120{1'b1}},194'b0};
  10'd589: road_rom_data = {199'b0,{120{1'b1}},193'b0};
  10'd590: road_rom_data = {199'b0,{120{1'b1}},193'b0};
  10'd591: road_rom_data = {200'b0,{120{1'b1}},192'b0};
  10'd592: road_rom_data = {201'b0,{120{1'b1}},191'b0};
  10'd593: road_rom_data = {202'b0,{120{1'b1}},190'b0};
  10'd594: road_rom_data = {202'b0,{120{1'b1}},190'b0};
  10'd595: road_rom_data = {203'b0,{120{1'b1}},189'b0};
  10'd596: road_rom_data = {204'b0,{120{1'b1}},188'b0};
  10'd597: road_rom_data = {205'b0,{120{1'b1}},187'b0};
  10'd598: road_rom_data = {205'b0,{120{1'b1}},187'b0};
  10'd599: road_rom_data = {206'b0,{120{1'b1}},186'b0};
  10'd600: road_rom_data = {207'b0,{120{1'b1}},185'b0};
  10'd601: road_rom_data = {208'b0,{120{1'b1}},184'b0};
  10'd602: road_rom_data = {208'b0,{120{1'b1}},184'b0};
  10'd603: road_rom_data = {209'b0,{120{1'b1}},183'b0};
  10'd604: road_rom_data = {210'b0,{120{1'b1}},182'b0};
  10'd605: road_rom_data = {211'b0,{120{1'b1}},181'b0};
  10'd606: road_rom_data = {211'b0,{120{1'b1}},181'b0};
  10'd607: road_rom_data = {212'b0,{120{1'b1}},180'b0};
  10'd608: road_rom_data = {213'b0,{120{1'b1}},179'b0};
  10'd609: road_rom_data = {214'b0,{120{1'b1}},178'b0};
  10'd610: road_rom_data = {214'b0,{120{1'b1}},178'b0};
  10'd611: road_rom_data = {215'b0,{120{1'b1}},177'b0};
  10'd612: road_rom_data = {216'b0,{120{1'b1}},176'b0};
  10'd613: road_rom_data = {216'b0,{120{1'b1}},176'b0};
  10'd614: road_rom_data = {217'b0,{120{1'b1}},175'b0};
  10'd615: road_rom_data = {218'b0,{120{1'b1}},174'b0};
  10'd616: road_rom_data = {218'b0,{120{1'b1}},174'b0};
  10'd617: road_rom_data = {219'b0,{120{1'b1}},173'b0};
  10'd618: road_rom_data = {220'b0,{120{1'b1}},172'b0};
  10'd619: road_rom_data = {220'b0,{120{1'b1}},172'b0};
  10'd620: road_rom_data = {221'b0,{120{1'b1}},171'b0};
  10'd621: road_rom_data = {222'b0,{120{1'b1}},170'b0};
  10'd622: road_rom_data = {222'b0,{120{1'b1}},170'b0};
  10'd623: road_rom_data = {223'b0,{120{1'b1}},169'b0};
  10'd624: road_rom_data = {224'b0,{120{1'b1}},168'b0};
  10'd625: road_rom_data = {224'b0,{120{1'b1}},168'b0};
  10'd626: road_rom_data = {225'b0,{120{1'b1}},167'b0};
  10'd627: road_rom_data = {226'b0,{120{1'b1}},166'b0};
  10'd628: road_rom_data = {226'b0,{120{1'b1}},166'b0};
  10'd629: road_rom_data = {227'b0,{120{1'b1}},165'b0};
  10'd630: road_rom_data = {227'b0,{120{1'b1}},165'b0};
  10'd631: road_rom_data = {228'b0,{120{1'b1}},164'b0};
  10'd632: road_rom_data = {229'b0,{120{1'b1}},163'b0};
  10'd633: road_rom_data = {229'b0,{120{1'b1}},163'b0};
  10'd634: road_rom_data = {230'b0,{120{1'b1}},162'b0};
  10'd635: road_rom_data = {230'b0,{120{1'b1}},162'b0};
  10'd636: road_rom_data = {231'b0,{120{1'b1}},161'b0};
  10'd637: road_rom_data = {232'b0,{120{1'b1}},160'b0};
  10'd638: road_rom_data = {232'b0,{120{1'b1}},160'b0};
  10'd639: road_rom_data = {233'b0,{120{1'b1}},159'b0};
  10'd640: road_rom_data = {233'b0,{120{1'b1}},159'b0};
  10'd641: road_rom_data = {234'b0,{120{1'b1}},158'b0};
  10'd642: road_rom_data = {234'b0,{120{1'b1}},158'b0};
  10'd643: road_rom_data = {235'b0,{120{1'b1}},157'b0};
  10'd644: road_rom_data = {235'b0,{120{1'b1}},157'b0};
  10'd645: road_rom_data = {236'b0,{120{1'b1}},156'b0};
  10'd646: road_rom_data = {237'b0,{120{1'b1}},155'b0};
  10'd647: road_rom_data = {237'b0,{120{1'b1}},155'b0};
  10'd648: road_rom_data = {238'b0,{120{1'b1}},154'b0};
  10'd649: road_rom_data = {238'b0,{120{1'b1}},154'b0};
  10'd650: road_rom_data = {239'b0,{120{1'b1}},153'b0};
  10'd651: road_rom_data = {239'b0,{120{1'b1}},153'b0};
  10'd652: road_rom_data = {240'b0,{120{1'b1}},152'b0};
  10'd653: road_rom_data = {240'b0,{120{1'b1}},152'b0};
  10'd654: road_rom_data = {241'b0,{120{1'b1}},151'b0};
  10'd655: road_rom_data = {241'b0,{120{1'b1}},151'b0};
  10'd656: road_rom_data = {242'b0,{120{1'b1}},150'b0};
  10'd657: road_rom_data = {242'b0,{120{1'b1}},150'b0};
  10'd658: road_rom_data = {242'b0,{120{1'b1}},150'b0};
  10'd659: road_rom_data = {243'b0,{120{1'b1}},149'b0};
  10'd660: road_rom_data = {243'b0,{120{1'b1}},149'b0};
  10'd661: road_rom_data = {244'b0,{120{1'b1}},148'b0};
  10'd662: road_rom_data = {244'b0,{120{1'b1}},148'b0};
  10'd663: road_rom_data = {245'b0,{120{1'b1}},147'b0};
  10'd664: road_rom_data = {245'b0,{120{1'b1}},147'b0};
  10'd665: road_rom_data = {246'b0,{120{1'b1}},146'b0};
  10'd666: road_rom_data = {246'b0,{120{1'b1}},146'b0};
  10'd667: road_rom_data = {246'b0,{120{1'b1}},146'b0};
  10'd668: road_rom_data = {247'b0,{120{1'b1}},145'b0};
  10'd669: road_rom_data = {247'b0,{120{1'b1}},145'b0};
  10'd670: road_rom_data = {248'b0,{120{1'b1}},144'b0};
  10'd671: road_rom_data = {248'b0,{120{1'b1}},144'b0};
  10'd672: road_rom_data = {248'b0,{120{1'b1}},144'b0};
  10'd673: road_rom_data = {249'b0,{120{1'b1}},143'b0};
  10'd674: road_rom_data = {249'b0,{120{1'b1}},143'b0};
  10'd675: road_rom_data = {249'b0,{120{1'b1}},143'b0};
  10'd676: road_rom_data = {250'b0,{120{1'b1}},142'b0};
  10'd677: road_rom_data = {250'b0,{120{1'b1}},142'b0};
  10'd678: road_rom_data = {251'b0,{120{1'b1}},141'b0};
  10'd679: road_rom_data = {251'b0,{120{1'b1}},141'b0};
  10'd680: road_rom_data = {251'b0,{120{1'b1}},141'b0};
  10'd681: road_rom_data = {252'b0,{120{1'b1}},140'b0};
  10'd682: road_rom_data = {252'b0,{120{1'b1}},140'b0};
  10'd683: road_rom_data = {252'b0,{120{1'b1}},140'b0};
  10'd684: road_rom_data = {253'b0,{120{1'b1}},139'b0};
  10'd685: road_rom_data = {253'b0,{120{1'b1}},139'b0};
  10'd686: road_rom_data = {253'b0,{120{1'b1}},139'b0};
  10'd687: road_rom_data = {253'b0,{120{1'b1}},139'b0};
  10'd688: road_rom_data = {254'b0,{120{1'b1}},138'b0};
  10'd689: road_rom_data = {254'b0,{120{1'b1}},138'b0};
  10'd690: road_rom_data = {254'b0,{120{1'b1}},138'b0};
  10'd691: road_rom_data = {255'b0,{120{1'b1}},137'b0};
  10'd692: road_rom_data = {255'b0,{120{1'b1}},137'b0};
  10'd693: road_rom_data = {255'b0,{120{1'b1}},137'b0};
  10'd694: road_rom_data = {255'b0,{120{1'b1}},137'b0};
  10'd695: road_rom_data = {256'b0,{120{1'b1}},136'b0};
  10'd696: road_rom_data = {256'b0,{120{1'b1}},136'b0};
  10'd697: road_rom_data = {256'b0,{120{1'b1}},136'b0};
  10'd698: road_rom_data = {256'b0,{120{1'b1}},136'b0};
  10'd699: road_rom_data = {257'b0,{120{1'b1}},135'b0};
  10'd700: road_rom_data = {257'b0,{120{1'b1}},135'b0};
  10'd701: road_rom_data = {257'b0,{120{1'b1}},135'b0};
  10'd702: road_rom_data = {257'b0,{120{1'b1}},135'b0};
  10'd703: road_rom_data = {257'b0,{120{1'b1}},135'b0};
  10'd704: road_rom_data = {258'b0,{120{1'b1}},134'b0};
  10'd705: road_rom_data = {258'b0,{120{1'b1}},134'b0};
  10'd706: road_rom_data = {258'b0,{120{1'b1}},134'b0};
  10'd707: road_rom_data = {258'b0,{120{1'b1}},134'b0};
  10'd708: road_rom_data = {258'b0,{120{1'b1}},134'b0};
  10'd709: road_rom_data = {259'b0,{120{1'b1}},133'b0};
  10'd710: road_rom_data = {259'b0,{120{1'b1}},133'b0};
  10'd711: road_rom_data = {259'b0,{120{1'b1}},133'b0};
  10'd712: road_rom_data = {259'b0,{120{1'b1}},133'b0};
  10'd713: road_rom_data = {259'b0,{120{1'b1}},133'b0};
  10'd714: road_rom_data = {259'b0,{120{1'b1}},133'b0};
  10'd715: road_rom_data = {259'b0,{120{1'b1}},133'b0};
  10'd716: road_rom_data = {260'b0,{120{1'b1}},132'b0};
  10'd717: road_rom_data = {260'b0,{120{1'b1}},132'b0};
  10'd718: road_rom_data = {260'b0,{120{1'b1}},132'b0};
  10'd719: road_rom_data = {260'b0,{120{1'b1}},132'b0};
  10'd720: road_rom_data = {260'b0,{120{1'b1}},132'b0};
  10'd721: road_rom_data = {260'b0,{120{1'b1}},132'b0};
  10'd722: road_rom_data = {260'b0,{120{1'b1}},132'b0};
  10'd723: road_rom_data = {260'b0,{120{1'b1}},132'b0};
  10'd724: road_rom_data = {260'b0,{120{1'b1}},132'b0};
  10'd725: road_rom_data = {260'b0,{120{1'b1}},132'b0};
  10'd726: road_rom_data = {260'b0,{120{1'b1}},132'b0};
  10'd727: road_rom_data = {261'b0,{120{1'b1}},131'b0};
  10'd728: road_rom_data = {261'b0,{120{1'b1}},131'b0};
  10'd729: road_rom_data = {261'b0,{120{1'b1}},131'b0};
  10'd730: road_rom_data = {261'b0,{120{1'b1}},131'b0};
  10'd731: road_rom_data = {261'b0,{120{1'b1}},131'b0};
  10'd732: road_rom_data = {261'b0,{120{1'b1}},131'b0};
  10'd733: road_rom_data = {261'b0,{120{1'b1}},131'b0};
  10'd734: road_rom_data = {261'b0,{120{1'b1}},131'b0};
  10'd735: road_rom_data = {261'b0,{120{1'b1}},131'b0};
  10'd736: road_rom_data = {261'b0,{120{1'b1}},131'b0};
  10'd737: road_rom_data = {261'b0,{120{1'b1}},131'b0};
  10'd738: road_rom_data = {261'b0,{120{1'b1}},131'b0};
  10'd739: road_rom_data = {261'b0,{120{1'b1}},131'b0};
  10'd740: road_rom_data = {261'b0,{120{1'b1}},131'b0};
  10'd741: road_rom_data = {261'b0,{120{1'b1}},131'b0};
  10'd742: road_rom_data = {261'b0,{120{1'b1}},131'b0};
  10'd743: road_rom_data = {261'b0,{120{1'b1}},131'b0};
  10'd744: road_rom_data = {261'b0,{120{1'b1}},131'b0};
  10'd745: road_rom_data = {261'b0,{120{1'b1}},131'b0};
  10'd746: road_rom_data = {261'b0,{120{1'b1}},131'b0};
  10'd747: road_rom_data = {261'b0,{120{1'b1}},131'b0};
  10'd748: road_rom_data = {260'b0,{120{1'b1}},132'b0};
  10'd749: road_rom_data = {260'b0,{120{1'b1}},132'b0};
  10'd750: road_rom_data = {260'b0,{120{1'b1}},132'b0};
  10'd751: road_rom_data = {260'b0,{120{1'b1}},132'b0};
  10'd752: road_rom_data = {260'b0,{120{1'b1}},132'b0};
  10'd753: road_rom_data = {260'b0,{120{1'b1}},132'b0};
  10'd754: road_rom_data = {260'b0,{120{1'b1}},132'b0};
  10'd755: road_rom_data = {260'b0,{120{1'b1}},132'b0};
  10'd756: road_rom_data = {260'b0,{120{1'b1}},132'b0};
  10'd757: road_rom_data = {260'b0,{120{1'b1}},132'b0};
  10'd758: road_rom_data = {260'b0,{120{1'b1}},132'b0};
  10'd759: road_rom_data = {259'b0,{120{1'b1}},133'b0};
  10'd760: road_rom_data = {259'b0,{120{1'b1}},133'b0};
  10'd761: road_rom_data = {259'b0,{120{1'b1}},133'b0};
  10'd762: road_rom_data = {259'b0,{120{1'b1}},133'b0};
  10'd763: road_rom_data = {259'b0,{120{1'b1}},133'b0};
  10'd764: road_rom_data = {259'b0,{120{1'b1}},133'b0};
  10'd765: road_rom_data = {259'b0,{120{1'b1}},133'b0};
  10'd766: road_rom_data = {258'b0,{120{1'b1}},134'b0};
  10'd767: road_rom_data = {258'b0,{120{1'b1}},134'b0};
  10'd768: road_rom_data = {258'b0,{120{1'b1}},134'b0};
  10'd769: road_rom_data = {258'b0,{120{1'b1}},134'b0};
  10'd770: road_rom_data = {258'b0,{120{1'b1}},134'b0};
  10'd771: road_rom_data = {258'b0,{120{1'b1}},134'b0};
  10'd772: road_rom_data = {257'b0,{120{1'b1}},135'b0};
  10'd773: road_rom_data = {257'b0,{120{1'b1}},135'b0};
  10'd774: road_rom_data = {257'b0,{120{1'b1}},135'b0};
  10'd775: road_rom_data = {257'b0,{120{1'b1}},135'b0};
  10'd776: road_rom_data = {257'b0,{120{1'b1}},135'b0};
  10'd777: road_rom_data = {256'b0,{120{1'b1}},136'b0};
  10'd778: road_rom_data = {256'b0,{120{1'b1}},136'b0};
  10'd779: road_rom_data = {256'b0,{120{1'b1}},136'b0};
  10'd780: road_rom_data = {256'b0,{120{1'b1}},136'b0};
  10'd781: road_rom_data = {255'b0,{120{1'b1}},137'b0};
  10'd782: road_rom_data = {255'b0,{120{1'b1}},137'b0};
  10'd783: road_rom_data = {255'b0,{120{1'b1}},137'b0};
  10'd784: road_rom_data = {255'b0,{120{1'b1}},137'b0};
  10'd785: road_rom_data = {254'b0,{120{1'b1}},138'b0};
  10'd786: road_rom_data = {254'b0,{120{1'b1}},138'b0};
  10'd787: road_rom_data = {254'b0,{120{1'b1}},138'b0};
  10'd788: road_rom_data = {254'b0,{120{1'b1}},138'b0};
  10'd789: road_rom_data = {253'b0,{120{1'b1}},139'b0};
  10'd790: road_rom_data = {253'b0,{120{1'b1}},139'b0};
  10'd791: road_rom_data = {253'b0,{120{1'b1}},139'b0};
  10'd792: road_rom_data = {253'b0,{120{1'b1}},139'b0};
  10'd793: road_rom_data = {252'b0,{120{1'b1}},140'b0};
  10'd794: road_rom_data = {252'b0,{120{1'b1}},140'b0};
  10'd795: road_rom_data = {252'b0,{120{1'b1}},140'b0};
  10'd796: road_rom_data = {251'b0,{120{1'b1}},141'b0};
  10'd797: road_rom_data = {251'b0,{120{1'b1}},141'b0};
  10'd798: road_rom_data = {251'b0,{120{1'b1}},141'b0};
  10'd799: road_rom_data = {250'b0,{120{1'b1}},142'b0};
  10'd800: road_rom_data = {250'b0,{120{1'b1}},142'b0};
  10'd801: road_rom_data = {250'b0,{120{1'b1}},142'b0};
  10'd802: road_rom_data = {249'b0,{120{1'b1}},143'b0};
  10'd803: road_rom_data = {249'b0,{120{1'b1}},143'b0};
  10'd804: road_rom_data = {249'b0,{120{1'b1}},143'b0};
  10'd805: road_rom_data = {248'b0,{120{1'b1}},144'b0};
  10'd806: road_rom_data = {248'b0,{120{1'b1}},144'b0};
  10'd807: road_rom_data = {248'b0,{120{1'b1}},144'b0};
  10'd808: road_rom_data = {247'b0,{120{1'b1}},145'b0};
  10'd809: road_rom_data = {247'b0,{120{1'b1}},145'b0};
  10'd810: road_rom_data = {247'b0,{120{1'b1}},145'b0};
  10'd811: road_rom_data = {246'b0,{120{1'b1}},146'b0};
  10'd812: road_rom_data = {246'b0,{120{1'b1}},146'b0};
  10'd813: road_rom_data = {245'b0,{120{1'b1}},147'b0};
  10'd814: road_rom_data = {245'b0,{120{1'b1}},147'b0};
  10'd815: road_rom_data = {245'b0,{120{1'b1}},147'b0};
  10'd816: road_rom_data = {244'b0,{120{1'b1}},148'b0};
  10'd817: road_rom_data = {244'b0,{120{1'b1}},148'b0};
  10'd818: road_rom_data = {244'b0,{120{1'b1}},148'b0};
  10'd819: road_rom_data = {243'b0,{120{1'b1}},149'b0};
  10'd820: road_rom_data = {243'b0,{120{1'b1}},149'b0};
  10'd821: road_rom_data = {242'b0,{120{1'b1}},150'b0};
  10'd822: road_rom_data = {242'b0,{120{1'b1}},150'b0};
  10'd823: road_rom_data = {241'b0,{120{1'b1}},151'b0};
  10'd824: road_rom_data = {241'b0,{120{1'b1}},151'b0};
  10'd825: road_rom_data = {241'b0,{120{1'b1}},151'b0};
  10'd826: road_rom_data = {240'b0,{120{1'b1}},152'b0};
  10'd827: road_rom_data = {240'b0,{120{1'b1}},152'b0};
  10'd828: road_rom_data = {239'b0,{120{1'b1}},153'b0};
  10'd829: road_rom_data = {239'b0,{120{1'b1}},153'b0};
  10'd830: road_rom_data = {238'b0,{120{1'b1}},154'b0};
  10'd831: road_rom_data = {238'b0,{120{1'b1}},154'b0};
  10'd832: road_rom_data = {238'b0,{120{1'b1}},154'b0};
  10'd833: road_rom_data = {237'b0,{120{1'b1}},155'b0};
  10'd834: road_rom_data = {237'b0,{120{1'b1}},155'b0};
  10'd835: road_rom_data = {236'b0,{120{1'b1}},156'b0};
  10'd836: road_rom_data = {236'b0,{120{1'b1}},156'b0};
  10'd837: road_rom_data = {235'b0,{120{1'b1}},157'b0};
  10'd838: road_rom_data = {235'b0,{120{1'b1}},157'b0};
  10'd839: road_rom_data = {234'b0,{120{1'b1}},158'b0};
  10'd840: road_rom_data = {234'b0,{120{1'b1}},158'b0};
  10'd841: road_rom_data = {233'b0,{120{1'b1}},159'b0};
  10'd842: road_rom_data = {233'b0,{120{1'b1}},159'b0};
  10'd843: road_rom_data = {232'b0,{120{1'b1}},160'b0};
  10'd844: road_rom_data = {232'b0,{120{1'b1}},160'b0};
  10'd845: road_rom_data = {231'b0,{120{1'b1}},161'b0};
  10'd846: road_rom_data = {231'b0,{120{1'b1}},161'b0};
  10'd847: road_rom_data = {230'b0,{120{1'b1}},162'b0};
  10'd848: road_rom_data = {230'b0,{120{1'b1}},162'b0};
  10'd849: road_rom_data = {229'b0,{120{1'b1}},163'b0};
  10'd850: road_rom_data = {229'b0,{120{1'b1}},163'b0};
  10'd851: road_rom_data = {228'b0,{120{1'b1}},164'b0};
  10'd852: road_rom_data = {228'b0,{120{1'b1}},164'b0};
  10'd853: road_rom_data = {227'b0,{120{1'b1}},165'b0};
  10'd854: road_rom_data = {227'b0,{120{1'b1}},165'b0};
  10'd855: road_rom_data = {226'b0,{120{1'b1}},166'b0};
  10'd856: road_rom_data = {226'b0,{120{1'b1}},166'b0};
  10'd857: road_rom_data = {225'b0,{120{1'b1}},167'b0};
  10'd858: road_rom_data = {225'b0,{120{1'b1}},167'b0};
  10'd859: road_rom_data = {224'b0,{120{1'b1}},168'b0};
  10'd860: road_rom_data = {224'b0,{120{1'b1}},168'b0};
  10'd861: road_rom_data = {223'b0,{120{1'b1}},169'b0};
  10'd862: road_rom_data = {223'b0,{120{1'b1}},169'b0};
  10'd863: road_rom_data = {222'b0,{120{1'b1}},170'b0};
  10'd864: road_rom_data = {222'b0,{120{1'b1}},170'b0};
  10'd865: road_rom_data = {221'b0,{120{1'b1}},171'b0};
  10'd866: road_rom_data = {221'b0,{120{1'b1}},171'b0};
  10'd867: road_rom_data = {220'b0,{120{1'b1}},172'b0};
  10'd868: road_rom_data = {219'b0,{120{1'b1}},173'b0};
  10'd869: road_rom_data = {219'b0,{120{1'b1}},173'b0};
  10'd870: road_rom_data = {218'b0,{120{1'b1}},174'b0};
  10'd871: road_rom_data = {218'b0,{120{1'b1}},174'b0};
  10'd872: road_rom_data = {217'b0,{120{1'b1}},175'b0};
  10'd873: road_rom_data = {217'b0,{120{1'b1}},175'b0};
  10'd874: road_rom_data = {216'b0,{120{1'b1}},176'b0};
  10'd875: road_rom_data = {216'b0,{120{1'b1}},176'b0};
  10'd876: road_rom_data = {215'b0,{120{1'b1}},177'b0};
  10'd877: road_rom_data = {215'b0,{120{1'b1}},177'b0};
  10'd878: road_rom_data = {214'b0,{120{1'b1}},178'b0};
  10'd879: road_rom_data = {213'b0,{120{1'b1}},179'b0};
  10'd880: road_rom_data = {213'b0,{120{1'b1}},179'b0};
  10'd881: road_rom_data = {212'b0,{120{1'b1}},180'b0};
  10'd882: road_rom_data = {212'b0,{120{1'b1}},180'b0};
  10'd883: road_rom_data = {211'b0,{120{1'b1}},181'b0};
  10'd884: road_rom_data = {211'b0,{120{1'b1}},181'b0};
  10'd885: road_rom_data = {210'b0,{120{1'b1}},182'b0};
  10'd886: road_rom_data = {209'b0,{120{1'b1}},183'b0};
  10'd887: road_rom_data = {209'b0,{120{1'b1}},183'b0};
  10'd888: road_rom_data = {208'b0,{120{1'b1}},184'b0};
  10'd889: road_rom_data = {208'b0,{120{1'b1}},184'b0};
  10'd890: road_rom_data = {207'b0,{120{1'b1}},185'b0};
  10'd891: road_rom_data = {207'b0,{120{1'b1}},185'b0};
  10'd892: road_rom_data = {206'b0,{120{1'b1}},186'b0};
  10'd893: road_rom_data = {205'b0,{120{1'b1}},187'b0};
  10'd894: road_rom_data = {205'b0,{120{1'b1}},187'b0};
  10'd895: road_rom_data = {204'b0,{120{1'b1}},188'b0};
  10'd896: road_rom_data = {204'b0,{120{1'b1}},188'b0};
  10'd897: road_rom_data = {203'b0,{120{1'b1}},189'b0};
  10'd898: road_rom_data = {203'b0,{120{1'b1}},189'b0};
  10'd899: road_rom_data = {202'b0,{120{1'b1}},190'b0};
  10'd900: road_rom_data = {201'b0,{120{1'b1}},191'b0};
  10'd901: road_rom_data = {201'b0,{120{1'b1}},191'b0};
  10'd902: road_rom_data = {200'b0,{120{1'b1}},192'b0};
  10'd903: road_rom_data = {200'b0,{120{1'b1}},192'b0};
  10'd904: road_rom_data = {199'b0,{120{1'b1}},193'b0};
  10'd905: road_rom_data = {198'b0,{120{1'b1}},194'b0};
  10'd906: road_rom_data = {198'b0,{120{1'b1}},194'b0};
  10'd907: road_rom_data = {197'b0,{120{1'b1}},195'b0};
  10'd908: road_rom_data = {197'b0,{120{1'b1}},195'b0};
  10'd909: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd910: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd911: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd912: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd913: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd914: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd915: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd916: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd917: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd918: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd919: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd920: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd921: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd922: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd923: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd924: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd925: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd926: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd927: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd928: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd929: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd930: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd931: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd932: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd933: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd934: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd935: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd936: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd937: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd938: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd939: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd940: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd941: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd942: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd943: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd944: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd945: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd946: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd947: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd948: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd949: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd950: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd951: road_rom_data = {200'b0,{112{1'b1}},200'b0};
  10'd952: road_rom_data = {200'b0,{112{1'b1}},200'b0};
  10'd953: road_rom_data = {200'b0,{112{1'b1}},200'b0};
  10'd954: road_rom_data = {200'b0,{112{1'b1}},200'b0};
  10'd955: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd956: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd957: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd958: road_rom_data = {196'b0,{120{1'b1}},196'b0};
  10'd959: road_rom_data = {196'b0,{120{1'b1}},196'b0};
      default: road_rom_data = 512'b0; //no road
  endcase
  

endmodule
